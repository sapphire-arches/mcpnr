// IO modules
(* blackbox, keep *)
module MCPNR_SWITCHES (
  output wire [NSWITCH-1:0] O
);
  parameter POS_X = 0;
  parameter POS_Y = 0;
  parameter POS_Z = 0;
  parameter NSWITCH = 1;
endmodule

(* blackbox, keep *)
module MCPNR_LIGHTS (
  input wire [NLIGHT-1:0] I
);
  parameter POS_X = 0;
  parameter POS_Y = 0;
  parameter POS_Z = 0;
  parameter NLIGHT = 1;
endmodule

// Functional modules.
// The names of these modules should correspond exactly with structure files in
// ./structures
//
// It's best if the order matches the one in minecraft.lib
// TODO: these should be autogenerated from the liberty function expressions

(* lib_blackbox, keep *)
module \gate_not.nbt (
  input  wire A,
  output wire Y
);
`ifndef BLACKBOX
  assign A = !Y;
`endif
endmodule

(* lib_blackbox, keep *)
module \gate_nand_i2.nbt (
  input  wire A, B,
  output wire Y
);
`ifndef BLACKBOX
  assign Y = !(A & B);
`endif
endmodule

(* lib_blackbox, keep *)
module \gate_nor_i2.nbt (
  input  wire A, B,
  output wire Y
);
`ifndef BLACKBOX
  assign Y = !(A | B);
`endif
endmodule

(* lib_blackbox, keep *)
module \gate_xor.nbt (
  input  wire A, B,
  output wire Y
);
`ifndef BLACKBOX
  assign Y = A ^ B;
`endif
endmodule

(* abc9_flop, lib_whitebox *)
module \dff.nbt (
  input  wire C, D,
  output reg Q
);
  initial Q = 0;
  always @(posedge C)
    Q <= D;
endmodule

module test_adder (
  input  [7:0] A, B,
  output [8:0] Y
);
  assign Y = A + B;
endmodule
